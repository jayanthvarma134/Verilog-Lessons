// AND gate

module and_b(out, x, y);
    input x, y;
    output out;
    assign out = x & y;
endmodule
